magic
tech sky130A
magscale 1 2
timestamp 1654670577
<< obsli1 >>
rect 1104 2159 358892 317713
<< obsm1 >>
rect 290 1368 359614 317892
<< metal2 >>
rect 1582 319200 1638 320000
rect 4710 319200 4766 320000
rect 7838 319200 7894 320000
rect 10966 319200 11022 320000
rect 14186 319200 14242 320000
rect 17314 319200 17370 320000
rect 20442 319200 20498 320000
rect 23662 319200 23718 320000
rect 26790 319200 26846 320000
rect 29918 319200 29974 320000
rect 33138 319200 33194 320000
rect 36266 319200 36322 320000
rect 39394 319200 39450 320000
rect 42614 319200 42670 320000
rect 45742 319200 45798 320000
rect 48870 319200 48926 320000
rect 52090 319200 52146 320000
rect 55218 319200 55274 320000
rect 58346 319200 58402 320000
rect 61566 319200 61622 320000
rect 64694 319200 64750 320000
rect 67822 319200 67878 320000
rect 71042 319200 71098 320000
rect 74170 319200 74226 320000
rect 77298 319200 77354 320000
rect 80518 319200 80574 320000
rect 83646 319200 83702 320000
rect 86774 319200 86830 320000
rect 89994 319200 90050 320000
rect 93122 319200 93178 320000
rect 96250 319200 96306 320000
rect 99470 319200 99526 320000
rect 102598 319200 102654 320000
rect 105726 319200 105782 320000
rect 108946 319200 109002 320000
rect 112074 319200 112130 320000
rect 115202 319200 115258 320000
rect 118422 319200 118478 320000
rect 121550 319200 121606 320000
rect 124678 319200 124734 320000
rect 127806 319200 127862 320000
rect 131026 319200 131082 320000
rect 134154 319200 134210 320000
rect 137282 319200 137338 320000
rect 140502 319200 140558 320000
rect 143630 319200 143686 320000
rect 146758 319200 146814 320000
rect 149978 319200 150034 320000
rect 153106 319200 153162 320000
rect 156234 319200 156290 320000
rect 159454 319200 159510 320000
rect 162582 319200 162638 320000
rect 165710 319200 165766 320000
rect 168930 319200 168986 320000
rect 172058 319200 172114 320000
rect 175186 319200 175242 320000
rect 178406 319200 178462 320000
rect 181534 319200 181590 320000
rect 184662 319200 184718 320000
rect 187882 319200 187938 320000
rect 191010 319200 191066 320000
rect 194138 319200 194194 320000
rect 197358 319200 197414 320000
rect 200486 319200 200542 320000
rect 203614 319200 203670 320000
rect 206834 319200 206890 320000
rect 209962 319200 210018 320000
rect 213090 319200 213146 320000
rect 216310 319200 216366 320000
rect 219438 319200 219494 320000
rect 222566 319200 222622 320000
rect 225786 319200 225842 320000
rect 228914 319200 228970 320000
rect 232042 319200 232098 320000
rect 235262 319200 235318 320000
rect 238390 319200 238446 320000
rect 241518 319200 241574 320000
rect 244646 319200 244702 320000
rect 247866 319200 247922 320000
rect 250994 319200 251050 320000
rect 254122 319200 254178 320000
rect 257342 319200 257398 320000
rect 260470 319200 260526 320000
rect 263598 319200 263654 320000
rect 266818 319200 266874 320000
rect 269946 319200 270002 320000
rect 273074 319200 273130 320000
rect 276294 319200 276350 320000
rect 279422 319200 279478 320000
rect 282550 319200 282606 320000
rect 285770 319200 285826 320000
rect 288898 319200 288954 320000
rect 292026 319200 292082 320000
rect 295246 319200 295302 320000
rect 298374 319200 298430 320000
rect 301502 319200 301558 320000
rect 304722 319200 304778 320000
rect 307850 319200 307906 320000
rect 310978 319200 311034 320000
rect 314198 319200 314254 320000
rect 317326 319200 317382 320000
rect 320454 319200 320510 320000
rect 323674 319200 323730 320000
rect 326802 319200 326858 320000
rect 329930 319200 329986 320000
rect 333150 319200 333206 320000
rect 336278 319200 336334 320000
rect 339406 319200 339462 320000
rect 342626 319200 342682 320000
rect 345754 319200 345810 320000
rect 348882 319200 348938 320000
rect 352102 319200 352158 320000
rect 355230 319200 355286 320000
rect 358358 319200 358414 320000
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2410 0 2466 800
rect 3146 0 3202 800
rect 3882 0 3938 800
rect 4618 0 4674 800
rect 5354 0 5410 800
rect 6090 0 6146 800
rect 6826 0 6882 800
rect 7562 0 7618 800
rect 8298 0 8354 800
rect 9034 0 9090 800
rect 9770 0 9826 800
rect 10506 0 10562 800
rect 11242 0 11298 800
rect 11886 0 11942 800
rect 12622 0 12678 800
rect 13358 0 13414 800
rect 14094 0 14150 800
rect 14830 0 14886 800
rect 15566 0 15622 800
rect 16302 0 16358 800
rect 17038 0 17094 800
rect 17774 0 17830 800
rect 18510 0 18566 800
rect 19246 0 19302 800
rect 19982 0 20038 800
rect 20718 0 20774 800
rect 21454 0 21510 800
rect 22190 0 22246 800
rect 22926 0 22982 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25778 0 25834 800
rect 26514 0 26570 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31666 0 31722 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35990 0 36046 800
rect 36726 0 36782 800
rect 37462 0 37518 800
rect 38198 0 38254 800
rect 38934 0 38990 800
rect 39670 0 39726 800
rect 40406 0 40462 800
rect 41142 0 41198 800
rect 41878 0 41934 800
rect 42614 0 42670 800
rect 43350 0 43406 800
rect 44086 0 44142 800
rect 44822 0 44878 800
rect 45558 0 45614 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47674 0 47730 800
rect 48410 0 48466 800
rect 49146 0 49202 800
rect 49882 0 49938 800
rect 50618 0 50674 800
rect 51354 0 51410 800
rect 52090 0 52146 800
rect 52826 0 52882 800
rect 53562 0 53618 800
rect 54298 0 54354 800
rect 55034 0 55090 800
rect 55770 0 55826 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59358 0 59414 800
rect 60094 0 60150 800
rect 60830 0 60886 800
rect 61566 0 61622 800
rect 62302 0 62358 800
rect 63038 0 63094 800
rect 63774 0 63830 800
rect 64510 0 64566 800
rect 65246 0 65302 800
rect 65982 0 66038 800
rect 66718 0 66774 800
rect 67454 0 67510 800
rect 68190 0 68246 800
rect 68926 0 68982 800
rect 69662 0 69718 800
rect 70306 0 70362 800
rect 71042 0 71098 800
rect 71778 0 71834 800
rect 72514 0 72570 800
rect 73250 0 73306 800
rect 73986 0 74042 800
rect 74722 0 74778 800
rect 75458 0 75514 800
rect 76194 0 76250 800
rect 76930 0 76986 800
rect 77666 0 77722 800
rect 78402 0 78458 800
rect 79138 0 79194 800
rect 79874 0 79930 800
rect 80610 0 80666 800
rect 81346 0 81402 800
rect 81990 0 82046 800
rect 82726 0 82782 800
rect 83462 0 83518 800
rect 84198 0 84254 800
rect 84934 0 84990 800
rect 85670 0 85726 800
rect 86406 0 86462 800
rect 87142 0 87198 800
rect 87878 0 87934 800
rect 88614 0 88670 800
rect 89350 0 89406 800
rect 90086 0 90142 800
rect 90822 0 90878 800
rect 91558 0 91614 800
rect 92294 0 92350 800
rect 93030 0 93086 800
rect 93674 0 93730 800
rect 94410 0 94466 800
rect 95146 0 95202 800
rect 95882 0 95938 800
rect 96618 0 96674 800
rect 97354 0 97410 800
rect 98090 0 98146 800
rect 98826 0 98882 800
rect 99562 0 99618 800
rect 100298 0 100354 800
rect 101034 0 101090 800
rect 101770 0 101826 800
rect 102506 0 102562 800
rect 103242 0 103298 800
rect 103978 0 104034 800
rect 104714 0 104770 800
rect 105358 0 105414 800
rect 106094 0 106150 800
rect 106830 0 106886 800
rect 107566 0 107622 800
rect 108302 0 108358 800
rect 109038 0 109094 800
rect 109774 0 109830 800
rect 110510 0 110566 800
rect 111246 0 111302 800
rect 111982 0 112038 800
rect 112718 0 112774 800
rect 113454 0 113510 800
rect 114190 0 114246 800
rect 114926 0 114982 800
rect 115662 0 115718 800
rect 116398 0 116454 800
rect 117042 0 117098 800
rect 117778 0 117834 800
rect 118514 0 118570 800
rect 119250 0 119306 800
rect 119986 0 120042 800
rect 120722 0 120778 800
rect 121458 0 121514 800
rect 122194 0 122250 800
rect 122930 0 122986 800
rect 123666 0 123722 800
rect 124402 0 124458 800
rect 125138 0 125194 800
rect 125874 0 125930 800
rect 126610 0 126666 800
rect 127346 0 127402 800
rect 127990 0 128046 800
rect 128726 0 128782 800
rect 129462 0 129518 800
rect 130198 0 130254 800
rect 130934 0 130990 800
rect 131670 0 131726 800
rect 132406 0 132462 800
rect 133142 0 133198 800
rect 133878 0 133934 800
rect 134614 0 134670 800
rect 135350 0 135406 800
rect 136086 0 136142 800
rect 136822 0 136878 800
rect 137558 0 137614 800
rect 138294 0 138350 800
rect 139030 0 139086 800
rect 139674 0 139730 800
rect 140410 0 140466 800
rect 141146 0 141202 800
rect 141882 0 141938 800
rect 142618 0 142674 800
rect 143354 0 143410 800
rect 144090 0 144146 800
rect 144826 0 144882 800
rect 145562 0 145618 800
rect 146298 0 146354 800
rect 147034 0 147090 800
rect 147770 0 147826 800
rect 148506 0 148562 800
rect 149242 0 149298 800
rect 149978 0 150034 800
rect 150714 0 150770 800
rect 151358 0 151414 800
rect 152094 0 152150 800
rect 152830 0 152886 800
rect 153566 0 153622 800
rect 154302 0 154358 800
rect 155038 0 155094 800
rect 155774 0 155830 800
rect 156510 0 156566 800
rect 157246 0 157302 800
rect 157982 0 158038 800
rect 158718 0 158774 800
rect 159454 0 159510 800
rect 160190 0 160246 800
rect 160926 0 160982 800
rect 161662 0 161718 800
rect 162398 0 162454 800
rect 163042 0 163098 800
rect 163778 0 163834 800
rect 164514 0 164570 800
rect 165250 0 165306 800
rect 165986 0 166042 800
rect 166722 0 166778 800
rect 167458 0 167514 800
rect 168194 0 168250 800
rect 168930 0 168986 800
rect 169666 0 169722 800
rect 170402 0 170458 800
rect 171138 0 171194 800
rect 171874 0 171930 800
rect 172610 0 172666 800
rect 173346 0 173402 800
rect 174082 0 174138 800
rect 174726 0 174782 800
rect 175462 0 175518 800
rect 176198 0 176254 800
rect 176934 0 176990 800
rect 177670 0 177726 800
rect 178406 0 178462 800
rect 179142 0 179198 800
rect 179878 0 179934 800
rect 180614 0 180670 800
rect 181350 0 181406 800
rect 182086 0 182142 800
rect 182822 0 182878 800
rect 183558 0 183614 800
rect 184294 0 184350 800
rect 185030 0 185086 800
rect 185766 0 185822 800
rect 186410 0 186466 800
rect 187146 0 187202 800
rect 187882 0 187938 800
rect 188618 0 188674 800
rect 189354 0 189410 800
rect 190090 0 190146 800
rect 190826 0 190882 800
rect 191562 0 191618 800
rect 192298 0 192354 800
rect 193034 0 193090 800
rect 193770 0 193826 800
rect 194506 0 194562 800
rect 195242 0 195298 800
rect 195978 0 196034 800
rect 196714 0 196770 800
rect 197450 0 197506 800
rect 198094 0 198150 800
rect 198830 0 198886 800
rect 199566 0 199622 800
rect 200302 0 200358 800
rect 201038 0 201094 800
rect 201774 0 201830 800
rect 202510 0 202566 800
rect 203246 0 203302 800
rect 203982 0 204038 800
rect 204718 0 204774 800
rect 205454 0 205510 800
rect 206190 0 206246 800
rect 206926 0 206982 800
rect 207662 0 207718 800
rect 208398 0 208454 800
rect 209134 0 209190 800
rect 209778 0 209834 800
rect 210514 0 210570 800
rect 211250 0 211306 800
rect 211986 0 212042 800
rect 212722 0 212778 800
rect 213458 0 213514 800
rect 214194 0 214250 800
rect 214930 0 214986 800
rect 215666 0 215722 800
rect 216402 0 216458 800
rect 217138 0 217194 800
rect 217874 0 217930 800
rect 218610 0 218666 800
rect 219346 0 219402 800
rect 220082 0 220138 800
rect 220818 0 220874 800
rect 221462 0 221518 800
rect 222198 0 222254 800
rect 222934 0 222990 800
rect 223670 0 223726 800
rect 224406 0 224462 800
rect 225142 0 225198 800
rect 225878 0 225934 800
rect 226614 0 226670 800
rect 227350 0 227406 800
rect 228086 0 228142 800
rect 228822 0 228878 800
rect 229558 0 229614 800
rect 230294 0 230350 800
rect 231030 0 231086 800
rect 231766 0 231822 800
rect 232502 0 232558 800
rect 233146 0 233202 800
rect 233882 0 233938 800
rect 234618 0 234674 800
rect 235354 0 235410 800
rect 236090 0 236146 800
rect 236826 0 236882 800
rect 237562 0 237618 800
rect 238298 0 238354 800
rect 239034 0 239090 800
rect 239770 0 239826 800
rect 240506 0 240562 800
rect 241242 0 241298 800
rect 241978 0 242034 800
rect 242714 0 242770 800
rect 243450 0 243506 800
rect 244094 0 244150 800
rect 244830 0 244886 800
rect 245566 0 245622 800
rect 246302 0 246358 800
rect 247038 0 247094 800
rect 247774 0 247830 800
rect 248510 0 248566 800
rect 249246 0 249302 800
rect 249982 0 250038 800
rect 250718 0 250774 800
rect 251454 0 251510 800
rect 252190 0 252246 800
rect 252926 0 252982 800
rect 253662 0 253718 800
rect 254398 0 254454 800
rect 255134 0 255190 800
rect 255778 0 255834 800
rect 256514 0 256570 800
rect 257250 0 257306 800
rect 257986 0 258042 800
rect 258722 0 258778 800
rect 259458 0 259514 800
rect 260194 0 260250 800
rect 260930 0 260986 800
rect 261666 0 261722 800
rect 262402 0 262458 800
rect 263138 0 263194 800
rect 263874 0 263930 800
rect 264610 0 264666 800
rect 265346 0 265402 800
rect 266082 0 266138 800
rect 266818 0 266874 800
rect 267462 0 267518 800
rect 268198 0 268254 800
rect 268934 0 268990 800
rect 269670 0 269726 800
rect 270406 0 270462 800
rect 271142 0 271198 800
rect 271878 0 271934 800
rect 272614 0 272670 800
rect 273350 0 273406 800
rect 274086 0 274142 800
rect 274822 0 274878 800
rect 275558 0 275614 800
rect 276294 0 276350 800
rect 277030 0 277086 800
rect 277766 0 277822 800
rect 278502 0 278558 800
rect 279146 0 279202 800
rect 279882 0 279938 800
rect 280618 0 280674 800
rect 281354 0 281410 800
rect 282090 0 282146 800
rect 282826 0 282882 800
rect 283562 0 283618 800
rect 284298 0 284354 800
rect 285034 0 285090 800
rect 285770 0 285826 800
rect 286506 0 286562 800
rect 287242 0 287298 800
rect 287978 0 288034 800
rect 288714 0 288770 800
rect 289450 0 289506 800
rect 290186 0 290242 800
rect 290830 0 290886 800
rect 291566 0 291622 800
rect 292302 0 292358 800
rect 293038 0 293094 800
rect 293774 0 293830 800
rect 294510 0 294566 800
rect 295246 0 295302 800
rect 295982 0 296038 800
rect 296718 0 296774 800
rect 297454 0 297510 800
rect 298190 0 298246 800
rect 298926 0 298982 800
rect 299662 0 299718 800
rect 300398 0 300454 800
rect 301134 0 301190 800
rect 301870 0 301926 800
rect 302514 0 302570 800
rect 303250 0 303306 800
rect 303986 0 304042 800
rect 304722 0 304778 800
rect 305458 0 305514 800
rect 306194 0 306250 800
rect 306930 0 306986 800
rect 307666 0 307722 800
rect 308402 0 308458 800
rect 309138 0 309194 800
rect 309874 0 309930 800
rect 310610 0 310666 800
rect 311346 0 311402 800
rect 312082 0 312138 800
rect 312818 0 312874 800
rect 313554 0 313610 800
rect 314198 0 314254 800
rect 314934 0 314990 800
rect 315670 0 315726 800
rect 316406 0 316462 800
rect 317142 0 317198 800
rect 317878 0 317934 800
rect 318614 0 318670 800
rect 319350 0 319406 800
rect 320086 0 320142 800
rect 320822 0 320878 800
rect 321558 0 321614 800
rect 322294 0 322350 800
rect 323030 0 323086 800
rect 323766 0 323822 800
rect 324502 0 324558 800
rect 325238 0 325294 800
rect 325882 0 325938 800
rect 326618 0 326674 800
rect 327354 0 327410 800
rect 328090 0 328146 800
rect 328826 0 328882 800
rect 329562 0 329618 800
rect 330298 0 330354 800
rect 331034 0 331090 800
rect 331770 0 331826 800
rect 332506 0 332562 800
rect 333242 0 333298 800
rect 333978 0 334034 800
rect 334714 0 334770 800
rect 335450 0 335506 800
rect 336186 0 336242 800
rect 336922 0 336978 800
rect 337566 0 337622 800
rect 338302 0 338358 800
rect 339038 0 339094 800
rect 339774 0 339830 800
rect 340510 0 340566 800
rect 341246 0 341302 800
rect 341982 0 342038 800
rect 342718 0 342774 800
rect 343454 0 343510 800
rect 344190 0 344246 800
rect 344926 0 344982 800
rect 345662 0 345718 800
rect 346398 0 346454 800
rect 347134 0 347190 800
rect 347870 0 347926 800
rect 348606 0 348662 800
rect 349250 0 349306 800
rect 349986 0 350042 800
rect 350722 0 350778 800
rect 351458 0 351514 800
rect 352194 0 352250 800
rect 352930 0 352986 800
rect 353666 0 353722 800
rect 354402 0 354458 800
rect 355138 0 355194 800
rect 355874 0 355930 800
rect 356610 0 356666 800
rect 357346 0 357402 800
rect 358082 0 358138 800
rect 358818 0 358874 800
rect 359554 0 359610 800
<< obsm2 >>
rect 296 319144 1526 319200
rect 1694 319144 4654 319200
rect 4822 319144 7782 319200
rect 7950 319144 10910 319200
rect 11078 319144 14130 319200
rect 14298 319144 17258 319200
rect 17426 319144 20386 319200
rect 20554 319144 23606 319200
rect 23774 319144 26734 319200
rect 26902 319144 29862 319200
rect 30030 319144 33082 319200
rect 33250 319144 36210 319200
rect 36378 319144 39338 319200
rect 39506 319144 42558 319200
rect 42726 319144 45686 319200
rect 45854 319144 48814 319200
rect 48982 319144 52034 319200
rect 52202 319144 55162 319200
rect 55330 319144 58290 319200
rect 58458 319144 61510 319200
rect 61678 319144 64638 319200
rect 64806 319144 67766 319200
rect 67934 319144 70986 319200
rect 71154 319144 74114 319200
rect 74282 319144 77242 319200
rect 77410 319144 80462 319200
rect 80630 319144 83590 319200
rect 83758 319144 86718 319200
rect 86886 319144 89938 319200
rect 90106 319144 93066 319200
rect 93234 319144 96194 319200
rect 96362 319144 99414 319200
rect 99582 319144 102542 319200
rect 102710 319144 105670 319200
rect 105838 319144 108890 319200
rect 109058 319144 112018 319200
rect 112186 319144 115146 319200
rect 115314 319144 118366 319200
rect 118534 319144 121494 319200
rect 121662 319144 124622 319200
rect 124790 319144 127750 319200
rect 127918 319144 130970 319200
rect 131138 319144 134098 319200
rect 134266 319144 137226 319200
rect 137394 319144 140446 319200
rect 140614 319144 143574 319200
rect 143742 319144 146702 319200
rect 146870 319144 149922 319200
rect 150090 319144 153050 319200
rect 153218 319144 156178 319200
rect 156346 319144 159398 319200
rect 159566 319144 162526 319200
rect 162694 319144 165654 319200
rect 165822 319144 168874 319200
rect 169042 319144 172002 319200
rect 172170 319144 175130 319200
rect 175298 319144 178350 319200
rect 178518 319144 181478 319200
rect 181646 319144 184606 319200
rect 184774 319144 187826 319200
rect 187994 319144 190954 319200
rect 191122 319144 194082 319200
rect 194250 319144 197302 319200
rect 197470 319144 200430 319200
rect 200598 319144 203558 319200
rect 203726 319144 206778 319200
rect 206946 319144 209906 319200
rect 210074 319144 213034 319200
rect 213202 319144 216254 319200
rect 216422 319144 219382 319200
rect 219550 319144 222510 319200
rect 222678 319144 225730 319200
rect 225898 319144 228858 319200
rect 229026 319144 231986 319200
rect 232154 319144 235206 319200
rect 235374 319144 238334 319200
rect 238502 319144 241462 319200
rect 241630 319144 244590 319200
rect 244758 319144 247810 319200
rect 247978 319144 250938 319200
rect 251106 319144 254066 319200
rect 254234 319144 257286 319200
rect 257454 319144 260414 319200
rect 260582 319144 263542 319200
rect 263710 319144 266762 319200
rect 266930 319144 269890 319200
rect 270058 319144 273018 319200
rect 273186 319144 276238 319200
rect 276406 319144 279366 319200
rect 279534 319144 282494 319200
rect 282662 319144 285714 319200
rect 285882 319144 288842 319200
rect 289010 319144 291970 319200
rect 292138 319144 295190 319200
rect 295358 319144 298318 319200
rect 298486 319144 301446 319200
rect 301614 319144 304666 319200
rect 304834 319144 307794 319200
rect 307962 319144 310922 319200
rect 311090 319144 314142 319200
rect 314310 319144 317270 319200
rect 317438 319144 320398 319200
rect 320566 319144 323618 319200
rect 323786 319144 326746 319200
rect 326914 319144 329874 319200
rect 330042 319144 333094 319200
rect 333262 319144 336222 319200
rect 336390 319144 339350 319200
rect 339518 319144 342570 319200
rect 342738 319144 345698 319200
rect 345866 319144 348826 319200
rect 348994 319144 352046 319200
rect 352214 319144 355174 319200
rect 355342 319144 358302 319200
rect 358470 319144 359608 319200
rect 296 856 359608 319144
rect 406 734 882 856
rect 1050 734 1618 856
rect 1786 734 2354 856
rect 2522 734 3090 856
rect 3258 734 3826 856
rect 3994 734 4562 856
rect 4730 734 5298 856
rect 5466 734 6034 856
rect 6202 734 6770 856
rect 6938 734 7506 856
rect 7674 734 8242 856
rect 8410 734 8978 856
rect 9146 734 9714 856
rect 9882 734 10450 856
rect 10618 734 11186 856
rect 11354 734 11830 856
rect 11998 734 12566 856
rect 12734 734 13302 856
rect 13470 734 14038 856
rect 14206 734 14774 856
rect 14942 734 15510 856
rect 15678 734 16246 856
rect 16414 734 16982 856
rect 17150 734 17718 856
rect 17886 734 18454 856
rect 18622 734 19190 856
rect 19358 734 19926 856
rect 20094 734 20662 856
rect 20830 734 21398 856
rect 21566 734 22134 856
rect 22302 734 22870 856
rect 23038 734 23514 856
rect 23682 734 24250 856
rect 24418 734 24986 856
rect 25154 734 25722 856
rect 25890 734 26458 856
rect 26626 734 27194 856
rect 27362 734 27930 856
rect 28098 734 28666 856
rect 28834 734 29402 856
rect 29570 734 30138 856
rect 30306 734 30874 856
rect 31042 734 31610 856
rect 31778 734 32346 856
rect 32514 734 33082 856
rect 33250 734 33818 856
rect 33986 734 34554 856
rect 34722 734 35198 856
rect 35366 734 35934 856
rect 36102 734 36670 856
rect 36838 734 37406 856
rect 37574 734 38142 856
rect 38310 734 38878 856
rect 39046 734 39614 856
rect 39782 734 40350 856
rect 40518 734 41086 856
rect 41254 734 41822 856
rect 41990 734 42558 856
rect 42726 734 43294 856
rect 43462 734 44030 856
rect 44198 734 44766 856
rect 44934 734 45502 856
rect 45670 734 46238 856
rect 46406 734 46882 856
rect 47050 734 47618 856
rect 47786 734 48354 856
rect 48522 734 49090 856
rect 49258 734 49826 856
rect 49994 734 50562 856
rect 50730 734 51298 856
rect 51466 734 52034 856
rect 52202 734 52770 856
rect 52938 734 53506 856
rect 53674 734 54242 856
rect 54410 734 54978 856
rect 55146 734 55714 856
rect 55882 734 56450 856
rect 56618 734 57186 856
rect 57354 734 57922 856
rect 58090 734 58566 856
rect 58734 734 59302 856
rect 59470 734 60038 856
rect 60206 734 60774 856
rect 60942 734 61510 856
rect 61678 734 62246 856
rect 62414 734 62982 856
rect 63150 734 63718 856
rect 63886 734 64454 856
rect 64622 734 65190 856
rect 65358 734 65926 856
rect 66094 734 66662 856
rect 66830 734 67398 856
rect 67566 734 68134 856
rect 68302 734 68870 856
rect 69038 734 69606 856
rect 69774 734 70250 856
rect 70418 734 70986 856
rect 71154 734 71722 856
rect 71890 734 72458 856
rect 72626 734 73194 856
rect 73362 734 73930 856
rect 74098 734 74666 856
rect 74834 734 75402 856
rect 75570 734 76138 856
rect 76306 734 76874 856
rect 77042 734 77610 856
rect 77778 734 78346 856
rect 78514 734 79082 856
rect 79250 734 79818 856
rect 79986 734 80554 856
rect 80722 734 81290 856
rect 81458 734 81934 856
rect 82102 734 82670 856
rect 82838 734 83406 856
rect 83574 734 84142 856
rect 84310 734 84878 856
rect 85046 734 85614 856
rect 85782 734 86350 856
rect 86518 734 87086 856
rect 87254 734 87822 856
rect 87990 734 88558 856
rect 88726 734 89294 856
rect 89462 734 90030 856
rect 90198 734 90766 856
rect 90934 734 91502 856
rect 91670 734 92238 856
rect 92406 734 92974 856
rect 93142 734 93618 856
rect 93786 734 94354 856
rect 94522 734 95090 856
rect 95258 734 95826 856
rect 95994 734 96562 856
rect 96730 734 97298 856
rect 97466 734 98034 856
rect 98202 734 98770 856
rect 98938 734 99506 856
rect 99674 734 100242 856
rect 100410 734 100978 856
rect 101146 734 101714 856
rect 101882 734 102450 856
rect 102618 734 103186 856
rect 103354 734 103922 856
rect 104090 734 104658 856
rect 104826 734 105302 856
rect 105470 734 106038 856
rect 106206 734 106774 856
rect 106942 734 107510 856
rect 107678 734 108246 856
rect 108414 734 108982 856
rect 109150 734 109718 856
rect 109886 734 110454 856
rect 110622 734 111190 856
rect 111358 734 111926 856
rect 112094 734 112662 856
rect 112830 734 113398 856
rect 113566 734 114134 856
rect 114302 734 114870 856
rect 115038 734 115606 856
rect 115774 734 116342 856
rect 116510 734 116986 856
rect 117154 734 117722 856
rect 117890 734 118458 856
rect 118626 734 119194 856
rect 119362 734 119930 856
rect 120098 734 120666 856
rect 120834 734 121402 856
rect 121570 734 122138 856
rect 122306 734 122874 856
rect 123042 734 123610 856
rect 123778 734 124346 856
rect 124514 734 125082 856
rect 125250 734 125818 856
rect 125986 734 126554 856
rect 126722 734 127290 856
rect 127458 734 127934 856
rect 128102 734 128670 856
rect 128838 734 129406 856
rect 129574 734 130142 856
rect 130310 734 130878 856
rect 131046 734 131614 856
rect 131782 734 132350 856
rect 132518 734 133086 856
rect 133254 734 133822 856
rect 133990 734 134558 856
rect 134726 734 135294 856
rect 135462 734 136030 856
rect 136198 734 136766 856
rect 136934 734 137502 856
rect 137670 734 138238 856
rect 138406 734 138974 856
rect 139142 734 139618 856
rect 139786 734 140354 856
rect 140522 734 141090 856
rect 141258 734 141826 856
rect 141994 734 142562 856
rect 142730 734 143298 856
rect 143466 734 144034 856
rect 144202 734 144770 856
rect 144938 734 145506 856
rect 145674 734 146242 856
rect 146410 734 146978 856
rect 147146 734 147714 856
rect 147882 734 148450 856
rect 148618 734 149186 856
rect 149354 734 149922 856
rect 150090 734 150658 856
rect 150826 734 151302 856
rect 151470 734 152038 856
rect 152206 734 152774 856
rect 152942 734 153510 856
rect 153678 734 154246 856
rect 154414 734 154982 856
rect 155150 734 155718 856
rect 155886 734 156454 856
rect 156622 734 157190 856
rect 157358 734 157926 856
rect 158094 734 158662 856
rect 158830 734 159398 856
rect 159566 734 160134 856
rect 160302 734 160870 856
rect 161038 734 161606 856
rect 161774 734 162342 856
rect 162510 734 162986 856
rect 163154 734 163722 856
rect 163890 734 164458 856
rect 164626 734 165194 856
rect 165362 734 165930 856
rect 166098 734 166666 856
rect 166834 734 167402 856
rect 167570 734 168138 856
rect 168306 734 168874 856
rect 169042 734 169610 856
rect 169778 734 170346 856
rect 170514 734 171082 856
rect 171250 734 171818 856
rect 171986 734 172554 856
rect 172722 734 173290 856
rect 173458 734 174026 856
rect 174194 734 174670 856
rect 174838 734 175406 856
rect 175574 734 176142 856
rect 176310 734 176878 856
rect 177046 734 177614 856
rect 177782 734 178350 856
rect 178518 734 179086 856
rect 179254 734 179822 856
rect 179990 734 180558 856
rect 180726 734 181294 856
rect 181462 734 182030 856
rect 182198 734 182766 856
rect 182934 734 183502 856
rect 183670 734 184238 856
rect 184406 734 184974 856
rect 185142 734 185710 856
rect 185878 734 186354 856
rect 186522 734 187090 856
rect 187258 734 187826 856
rect 187994 734 188562 856
rect 188730 734 189298 856
rect 189466 734 190034 856
rect 190202 734 190770 856
rect 190938 734 191506 856
rect 191674 734 192242 856
rect 192410 734 192978 856
rect 193146 734 193714 856
rect 193882 734 194450 856
rect 194618 734 195186 856
rect 195354 734 195922 856
rect 196090 734 196658 856
rect 196826 734 197394 856
rect 197562 734 198038 856
rect 198206 734 198774 856
rect 198942 734 199510 856
rect 199678 734 200246 856
rect 200414 734 200982 856
rect 201150 734 201718 856
rect 201886 734 202454 856
rect 202622 734 203190 856
rect 203358 734 203926 856
rect 204094 734 204662 856
rect 204830 734 205398 856
rect 205566 734 206134 856
rect 206302 734 206870 856
rect 207038 734 207606 856
rect 207774 734 208342 856
rect 208510 734 209078 856
rect 209246 734 209722 856
rect 209890 734 210458 856
rect 210626 734 211194 856
rect 211362 734 211930 856
rect 212098 734 212666 856
rect 212834 734 213402 856
rect 213570 734 214138 856
rect 214306 734 214874 856
rect 215042 734 215610 856
rect 215778 734 216346 856
rect 216514 734 217082 856
rect 217250 734 217818 856
rect 217986 734 218554 856
rect 218722 734 219290 856
rect 219458 734 220026 856
rect 220194 734 220762 856
rect 220930 734 221406 856
rect 221574 734 222142 856
rect 222310 734 222878 856
rect 223046 734 223614 856
rect 223782 734 224350 856
rect 224518 734 225086 856
rect 225254 734 225822 856
rect 225990 734 226558 856
rect 226726 734 227294 856
rect 227462 734 228030 856
rect 228198 734 228766 856
rect 228934 734 229502 856
rect 229670 734 230238 856
rect 230406 734 230974 856
rect 231142 734 231710 856
rect 231878 734 232446 856
rect 232614 734 233090 856
rect 233258 734 233826 856
rect 233994 734 234562 856
rect 234730 734 235298 856
rect 235466 734 236034 856
rect 236202 734 236770 856
rect 236938 734 237506 856
rect 237674 734 238242 856
rect 238410 734 238978 856
rect 239146 734 239714 856
rect 239882 734 240450 856
rect 240618 734 241186 856
rect 241354 734 241922 856
rect 242090 734 242658 856
rect 242826 734 243394 856
rect 243562 734 244038 856
rect 244206 734 244774 856
rect 244942 734 245510 856
rect 245678 734 246246 856
rect 246414 734 246982 856
rect 247150 734 247718 856
rect 247886 734 248454 856
rect 248622 734 249190 856
rect 249358 734 249926 856
rect 250094 734 250662 856
rect 250830 734 251398 856
rect 251566 734 252134 856
rect 252302 734 252870 856
rect 253038 734 253606 856
rect 253774 734 254342 856
rect 254510 734 255078 856
rect 255246 734 255722 856
rect 255890 734 256458 856
rect 256626 734 257194 856
rect 257362 734 257930 856
rect 258098 734 258666 856
rect 258834 734 259402 856
rect 259570 734 260138 856
rect 260306 734 260874 856
rect 261042 734 261610 856
rect 261778 734 262346 856
rect 262514 734 263082 856
rect 263250 734 263818 856
rect 263986 734 264554 856
rect 264722 734 265290 856
rect 265458 734 266026 856
rect 266194 734 266762 856
rect 266930 734 267406 856
rect 267574 734 268142 856
rect 268310 734 268878 856
rect 269046 734 269614 856
rect 269782 734 270350 856
rect 270518 734 271086 856
rect 271254 734 271822 856
rect 271990 734 272558 856
rect 272726 734 273294 856
rect 273462 734 274030 856
rect 274198 734 274766 856
rect 274934 734 275502 856
rect 275670 734 276238 856
rect 276406 734 276974 856
rect 277142 734 277710 856
rect 277878 734 278446 856
rect 278614 734 279090 856
rect 279258 734 279826 856
rect 279994 734 280562 856
rect 280730 734 281298 856
rect 281466 734 282034 856
rect 282202 734 282770 856
rect 282938 734 283506 856
rect 283674 734 284242 856
rect 284410 734 284978 856
rect 285146 734 285714 856
rect 285882 734 286450 856
rect 286618 734 287186 856
rect 287354 734 287922 856
rect 288090 734 288658 856
rect 288826 734 289394 856
rect 289562 734 290130 856
rect 290298 734 290774 856
rect 290942 734 291510 856
rect 291678 734 292246 856
rect 292414 734 292982 856
rect 293150 734 293718 856
rect 293886 734 294454 856
rect 294622 734 295190 856
rect 295358 734 295926 856
rect 296094 734 296662 856
rect 296830 734 297398 856
rect 297566 734 298134 856
rect 298302 734 298870 856
rect 299038 734 299606 856
rect 299774 734 300342 856
rect 300510 734 301078 856
rect 301246 734 301814 856
rect 301982 734 302458 856
rect 302626 734 303194 856
rect 303362 734 303930 856
rect 304098 734 304666 856
rect 304834 734 305402 856
rect 305570 734 306138 856
rect 306306 734 306874 856
rect 307042 734 307610 856
rect 307778 734 308346 856
rect 308514 734 309082 856
rect 309250 734 309818 856
rect 309986 734 310554 856
rect 310722 734 311290 856
rect 311458 734 312026 856
rect 312194 734 312762 856
rect 312930 734 313498 856
rect 313666 734 314142 856
rect 314310 734 314878 856
rect 315046 734 315614 856
rect 315782 734 316350 856
rect 316518 734 317086 856
rect 317254 734 317822 856
rect 317990 734 318558 856
rect 318726 734 319294 856
rect 319462 734 320030 856
rect 320198 734 320766 856
rect 320934 734 321502 856
rect 321670 734 322238 856
rect 322406 734 322974 856
rect 323142 734 323710 856
rect 323878 734 324446 856
rect 324614 734 325182 856
rect 325350 734 325826 856
rect 325994 734 326562 856
rect 326730 734 327298 856
rect 327466 734 328034 856
rect 328202 734 328770 856
rect 328938 734 329506 856
rect 329674 734 330242 856
rect 330410 734 330978 856
rect 331146 734 331714 856
rect 331882 734 332450 856
rect 332618 734 333186 856
rect 333354 734 333922 856
rect 334090 734 334658 856
rect 334826 734 335394 856
rect 335562 734 336130 856
rect 336298 734 336866 856
rect 337034 734 337510 856
rect 337678 734 338246 856
rect 338414 734 338982 856
rect 339150 734 339718 856
rect 339886 734 340454 856
rect 340622 734 341190 856
rect 341358 734 341926 856
rect 342094 734 342662 856
rect 342830 734 343398 856
rect 343566 734 344134 856
rect 344302 734 344870 856
rect 345038 734 345606 856
rect 345774 734 346342 856
rect 346510 734 347078 856
rect 347246 734 347814 856
rect 347982 734 348550 856
rect 348718 734 349194 856
rect 349362 734 349930 856
rect 350098 734 350666 856
rect 350834 734 351402 856
rect 351570 734 352138 856
rect 352306 734 352874 856
rect 353042 734 353610 856
rect 353778 734 354346 856
rect 354514 734 355082 856
rect 355250 734 355818 856
rect 355986 734 356554 856
rect 356722 734 357290 856
rect 357458 734 358026 856
rect 358194 734 358762 856
rect 358930 734 359498 856
<< obsm3 >>
rect 4210 2143 354526 317729
<< metal4 >>
rect 4208 2128 4528 317744
rect 14208 2128 14528 317744
rect 24208 2128 24528 317744
rect 34208 2128 34528 317744
rect 44208 2128 44528 317744
rect 54208 2128 54528 317744
rect 64208 2128 64528 317744
rect 74208 2128 74528 317744
rect 84208 2128 84528 317744
rect 94208 2128 94528 317744
rect 104208 2128 104528 317744
rect 114208 2128 114528 317744
rect 124208 2128 124528 317744
rect 134208 2128 134528 317744
rect 144208 2128 144528 317744
rect 154208 2128 154528 317744
rect 164208 2128 164528 317744
rect 174208 2128 174528 317744
rect 184208 2128 184528 317744
rect 194208 2128 194528 317744
rect 204208 2128 204528 317744
rect 214208 2128 214528 317744
rect 224208 2128 224528 317744
rect 234208 2128 234528 317744
rect 244208 2128 244528 317744
rect 254208 2128 254528 317744
rect 264208 2128 264528 317744
rect 274208 2128 274528 317744
rect 284208 2128 284528 317744
rect 294208 2128 294528 317744
rect 304208 2128 304528 317744
rect 314208 2128 314528 317744
rect 324208 2128 324528 317744
rect 334208 2128 334528 317744
rect 344208 2128 344528 317744
rect 354208 2128 354528 317744
<< obsm4 >>
rect 32995 31451 34128 302293
rect 34608 31451 44128 302293
rect 44608 31451 54128 302293
rect 54608 31451 64128 302293
rect 64608 31451 74128 302293
rect 74608 31451 84128 302293
rect 84608 31451 94128 302293
rect 94608 31451 104128 302293
rect 104608 31451 114128 302293
rect 114608 31451 124128 302293
rect 124608 31451 134128 302293
rect 134608 31451 144128 302293
rect 144608 31451 154128 302293
rect 154608 31451 164128 302293
rect 164608 31451 174128 302293
rect 174608 31451 184128 302293
rect 184608 31451 194128 302293
rect 194608 31451 204128 302293
rect 204608 31451 214128 302293
rect 214608 31451 224128 302293
rect 224608 31451 234128 302293
rect 234608 31451 244128 302293
rect 244608 31451 254128 302293
rect 254608 31451 264128 302293
rect 264608 31451 274128 302293
rect 274608 31451 284128 302293
rect 284608 31451 294128 302293
rect 294608 31451 304128 302293
rect 304608 31451 314128 302293
rect 314608 31451 324128 302293
rect 324608 31451 329485 302293
<< labels >>
rlabel metal2 s 1582 319200 1638 320000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 96250 319200 96306 320000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 105726 319200 105782 320000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 115202 319200 115258 320000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 124678 319200 124734 320000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 134154 319200 134210 320000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 143630 319200 143686 320000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 153106 319200 153162 320000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 162582 319200 162638 320000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 172058 319200 172114 320000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 181534 319200 181590 320000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 10966 319200 11022 320000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 191010 319200 191066 320000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 200486 319200 200542 320000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 209962 319200 210018 320000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 219438 319200 219494 320000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 228914 319200 228970 320000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 238390 319200 238446 320000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 247866 319200 247922 320000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 257342 319200 257398 320000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 266818 319200 266874 320000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 276294 319200 276350 320000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 20442 319200 20498 320000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 285770 319200 285826 320000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 295246 319200 295302 320000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 304722 319200 304778 320000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 314198 319200 314254 320000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 323674 319200 323730 320000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 333150 319200 333206 320000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 342626 319200 342682 320000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 352102 319200 352158 320000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 29918 319200 29974 320000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 39394 319200 39450 320000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 48870 319200 48926 320000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 58346 319200 58402 320000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 67822 319200 67878 320000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 77298 319200 77354 320000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 86774 319200 86830 320000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4710 319200 4766 320000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 99470 319200 99526 320000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 108946 319200 109002 320000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 118422 319200 118478 320000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 127806 319200 127862 320000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 137282 319200 137338 320000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 146758 319200 146814 320000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 156234 319200 156290 320000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 165710 319200 165766 320000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 175186 319200 175242 320000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 184662 319200 184718 320000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 14186 319200 14242 320000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 194138 319200 194194 320000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 203614 319200 203670 320000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 213090 319200 213146 320000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 222566 319200 222622 320000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 232042 319200 232098 320000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 241518 319200 241574 320000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 250994 319200 251050 320000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 260470 319200 260526 320000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 269946 319200 270002 320000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 279422 319200 279478 320000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 23662 319200 23718 320000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 288898 319200 288954 320000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 298374 319200 298430 320000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 307850 319200 307906 320000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 317326 319200 317382 320000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 326802 319200 326858 320000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 336278 319200 336334 320000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 345754 319200 345810 320000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 355230 319200 355286 320000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 33138 319200 33194 320000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 42614 319200 42670 320000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 52090 319200 52146 320000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 61566 319200 61622 320000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 71042 319200 71098 320000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 80518 319200 80574 320000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 89994 319200 90050 320000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 7838 319200 7894 320000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 102598 319200 102654 320000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 112074 319200 112130 320000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 121550 319200 121606 320000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 131026 319200 131082 320000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 140502 319200 140558 320000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 149978 319200 150034 320000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 159454 319200 159510 320000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 168930 319200 168986 320000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 178406 319200 178462 320000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 187882 319200 187938 320000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 17314 319200 17370 320000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 197358 319200 197414 320000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 206834 319200 206890 320000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 216310 319200 216366 320000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 225786 319200 225842 320000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 235262 319200 235318 320000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 244646 319200 244702 320000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 254122 319200 254178 320000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 263598 319200 263654 320000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 273074 319200 273130 320000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 282550 319200 282606 320000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 26790 319200 26846 320000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 292026 319200 292082 320000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 301502 319200 301558 320000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 310978 319200 311034 320000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 320454 319200 320510 320000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 329930 319200 329986 320000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 339406 319200 339462 320000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 348882 319200 348938 320000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 358358 319200 358414 320000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 36266 319200 36322 320000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 45742 319200 45798 320000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 55218 319200 55274 320000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 64694 319200 64750 320000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 74170 319200 74226 320000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 83646 319200 83702 320000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 93122 319200 93178 320000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 358082 0 358138 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 358818 0 358874 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 359554 0 359610 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 296718 0 296774 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 298926 0 298982 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 301134 0 301190 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 303250 0 303306 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 305458 0 305514 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 307666 0 307722 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 309874 0 309930 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 312082 0 312138 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 314198 0 314254 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 316406 0 316462 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 318614 0 318670 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 320822 0 320878 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 323030 0 323086 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 325238 0 325294 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 329562 0 329618 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 331770 0 331826 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 333978 0 334034 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 338302 0 338358 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 340510 0 340566 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 342718 0 342774 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 344926 0 344982 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 347134 0 347190 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 351458 0 351514 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 353666 0 353722 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 355874 0 355930 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 231030 0 231086 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 235354 0 235410 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 244094 0 244150 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 250718 0 250774 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 252926 0 252982 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 255134 0 255190 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 259458 0 259514 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 261666 0 261722 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 263874 0 263930 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 266082 0 266138 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 272614 0 272670 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 274822 0 274878 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 279146 0 279202 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 283562 0 283618 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 285770 0 285826 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 287978 0 288034 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 290186 0 290242 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 292302 0 292358 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 297454 0 297510 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 299662 0 299718 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 301870 0 301926 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 303986 0 304042 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 306194 0 306250 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 308402 0 308458 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 310610 0 310666 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 312818 0 312874 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 314934 0 314990 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 317142 0 317198 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 319350 0 319406 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 321558 0 321614 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 323766 0 323822 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 325882 0 325938 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 328090 0 328146 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 330298 0 330354 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 332506 0 332562 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 334714 0 334770 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 336922 0 336978 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 339038 0 339094 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 341246 0 341302 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 343454 0 343510 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 345662 0 345718 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 347870 0 347926 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 349986 0 350042 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 352194 0 352250 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 354402 0 354458 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 356610 0 356666 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 155038 0 155094 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 163778 0 163834 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 181350 0 181406 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 185766 0 185822 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 187882 0 187938 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 190090 0 190146 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 194506 0 194562 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 198830 0 198886 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 203246 0 203302 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 209778 0 209834 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 211986 0 212042 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 220818 0 220874 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 222934 0 222990 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 225142 0 225198 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 231766 0 231822 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 236090 0 236146 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 238298 0 238354 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 242714 0 242770 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 244830 0 244886 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 247038 0 247094 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 249246 0 249302 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 253662 0 253718 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 255778 0 255834 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 257986 0 258042 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 260194 0 260250 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 264610 0 264666 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 266818 0 266874 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 271142 0 271198 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 273350 0 273406 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 275558 0 275614 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 277766 0 277822 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 279882 0 279938 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 282090 0 282146 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 284298 0 284354 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 286506 0 286562 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 288714 0 288770 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 290830 0 290886 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 293038 0 293094 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 295246 0 295302 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 302514 0 302570 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 304722 0 304778 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 306930 0 306986 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 309138 0 309194 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 311346 0 311402 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 313554 0 313610 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 315670 0 315726 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 317878 0 317934 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 320086 0 320142 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 324502 0 324558 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 326618 0 326674 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 328826 0 328882 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 331034 0 331090 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 333242 0 333298 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 335450 0 335506 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 337566 0 337622 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 339774 0 339830 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 341982 0 342038 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 344190 0 344246 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 346398 0 346454 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 348606 0 348662 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 350722 0 350778 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 352930 0 352986 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 355138 0 355194 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 357346 0 357402 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 212722 0 212778 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 221462 0 221518 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 225878 0 225934 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 230294 0 230350 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 243450 0 243506 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 247774 0 247830 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 256514 0 256570 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 258722 0 258778 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 260930 0 260986 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 267462 0 267518 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 271878 0 271934 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 278502 0 278558 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 285034 0 285090 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 287242 0 287298 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 289450 0 289506 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 293774 0 293830 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 244208 2128 244528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 264208 2128 264528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 284208 2128 284528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 304208 2128 304528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 324208 2128 324528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 344208 2128 344528 317744 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 34208 2128 34528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 54208 2128 54528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 74208 2128 74528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 94208 2128 94528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 114208 2128 114528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 134208 2128 134528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 154208 2128 154528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 174208 2128 174528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 194208 2128 194528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 214208 2128 214528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234208 2128 234528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 254208 2128 254528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 274208 2128 274528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 294208 2128 294528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 314208 2128 314528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 334208 2128 334528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 354208 2128 354528 317744 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 360000 320000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 142330200
string GDS_FILE /home/recep_linux/Desktop/mpw6_aes_rng/mpw6_crypto_rng/openlane/user_proj_example/runs/user_proj_example/results/signoff/user_proj_example.magic.gds
string GDS_START 1342528
<< end >>

